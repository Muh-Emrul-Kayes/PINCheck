# 
# ******************************************************************************
# *                                                                            *
# *                   Copyright (C) 2004-2016, Nangate Inc.                    *
# *                           All rights reserved.                             *
# *                                                                            *
# * Nangate and the Nangate logo are trademarks of Nangate Inc.                *
# *                                                                            *
# * All trademarks, logos, software marks, and trade names (collectively the   *
# * "Marks") in this program are proprietary to Nangate or other respective    *
# * owners that have granted Nangate the right and license to use such Marks.  *
# * You are not permitted to use the Marks without the prior written consent   *
# * of Nangate or such third party that may own the Marks.                     *
# *                                                                            *
# * This file has been provided pursuant to a License Agreement containing     *
# * restrictions on its use. This file contains valuable trade secrets and     *
# * proprietary information of Nangate Inc., and is protected by U.S. and      *
# * international laws and/or treaties.                                        *
# *                                                                            *
# * The copyright notice(s) in this file does not indicate actual or intended  *
# * publication of this file.                                                  *
# *                                                                            *
# *       NGLibraryCreator, Development_version_64 - build 201509171155        *
# *                                                                            *
# ******************************************************************************
# 
# 
# Running on usdev01.nangate.us for user Guilherme Simoes Schlinker (gss).
# Local time is now Wed, 10 Feb 2016, 14:28:25.
# Main process id is 27110.

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO ISO_FENCE0N_X1_RVT_30
  CLASS core ;
  FOREIGN ISO_FENCE0N_X1_RVT_30 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CellTemplate ;
  SIZE 0.52 BY 0.8 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.00774 ;
    PORT
      LAYER M1 ;
        POLYGON 0.083 0.321 0.155 0.321 0.155 0.49 0.083 0.49  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.00774 ;
    PORT
      LAYER M1 ;
        POLYGON 0.207 0.323 0.273 0.323 0.273 0.49 0.207 0.49  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.040248 ;
    PORT
      LAYER M1 ;
        POLYGON 0.411 0.634 0.43 0.634 0.43 0.489 0.445 0.489 0.445 0.312 0.43 0.312 0.43 0.154 0.419 0.154 0.419 0.091 0.495 0.091 0.495 0.709 0.411 0.709  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 0.735 0.52 0.735 0.52 0.865 0 0.865  ;
      LAYER V1 ;
        POLYGON 0.04 0.775 0.09 0.775 0.09 0.825 0.04 0.825  ;
        POLYGON 0.17 0.775 0.22 0.775 0.22 0.825 0.17 0.825  ;
        POLYGON 0.3 0.775 0.35 0.775 0.35 0.825 0.3 0.825  ;
        POLYGON 0.43 0.775 0.48 0.775 0.48 0.825 0.43 0.825  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 -0.065 0.52 -0.065 0.52 0.065 0 0.065  ;
      LAYER V1 ;
        POLYGON 0.04 -0.025 0.09 -0.025 0.09 0.025 0.04 0.025  ;
        POLYGON 0.17 -0.025 0.22 -0.025 0.22 0.025 0.17 0.025  ;
        POLYGON 0.3 -0.025 0.35 -0.025 0.35 0.025 0.3 0.025  ;
        POLYGON 0.43 -0.025 0.48 -0.025 0.48 0.025 0.43 0.025  ;
    END
  END VSS
  OBS
      LAYER RVT ;
        POLYGON 0 0 0.52 0 0.52 0.8 0 0.8 ;
      LAYER M1 ;
        POLYGON 0.159 0.548 0.323 0.548 0.323 0.263 0.04 0.263 0.04 0.091 0.115 0.091 0.115 0.199 0.373 0.199 0.373 0.348 0.395 0.348 0.395 0.452 0.373 0.452 0.373 0.598 0.231 0.598 0.231 0.709 0.159 0.709  ;
        POLYGON 0 -0.033 0.52 -0.033 0.52 0.033 0.361 0.033 0.361 0.126 0.289 0.126 0.289 0.033 0 0.033  ;
        POLYGON 0 0.767 0.029 0.767 0.029 0.578 0.101 0.578 0.101 0.767 0.289 0.767 0.289 0.656 0.361 0.656 0.361 0.767 0.52 0.767 0.52 0.833 0 0.833  ;
  END
END ISO_FENCE0N_X1_RVT_30

MACRO ISO_FENCE0N_X2_RVT_30
  CLASS core ;
  FOREIGN ISO_FENCE0N_X2_RVT_30 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CellTemplate ;
  SIZE 0.65 BY 0.8 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.01548 ;
    PORT
      LAYER M1 ;
        POLYGON 0.083 0.321 0.155 0.321 0.155 0.483 0.083 0.483  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.01548 ;
    PORT
      LAYER M1 ;
        POLYGON 0.207 0.321 0.273 0.321 0.273 0.483 0.207 0.483  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.0516 ;
    PORT
      LAYER M1 ;
        POLYGON 0.423 0.475 0.556 0.475 0.556 0.269 0.423 0.269 0.423 0.091 0.489 0.091 0.489 0.219 0.606 0.219 0.606 0.525 0.489 0.525 0.489 0.709 0.423 0.709  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 0.735 0.65 0.735 0.65 0.865 0 0.865  ;
      LAYER V1 ;
        POLYGON 0.04 0.775 0.09 0.775 0.09 0.825 0.04 0.825  ;
        POLYGON 0.17 0.775 0.22 0.775 0.22 0.825 0.17 0.825  ;
        POLYGON 0.3 0.775 0.35 0.775 0.35 0.825 0.3 0.825  ;
        POLYGON 0.43 0.775 0.48 0.775 0.48 0.825 0.43 0.825  ;
        POLYGON 0.56 0.775 0.61 0.775 0.61 0.825 0.56 0.825  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 -0.065 0.65 -0.065 0.65 0.065 0 0.065  ;
      LAYER V1 ;
        POLYGON 0.04 -0.025 0.09 -0.025 0.09 0.025 0.04 0.025  ;
        POLYGON 0.17 -0.025 0.22 -0.025 0.22 0.025 0.17 0.025  ;
        POLYGON 0.3 -0.025 0.35 -0.025 0.35 0.025 0.3 0.025  ;
        POLYGON 0.43 -0.025 0.48 -0.025 0.48 0.025 0.43 0.025  ;
        POLYGON 0.56 -0.025 0.61 -0.025 0.61 0.025 0.56 0.025  ;
    END
  END VSS
  OBS
      LAYER RVT ;
        POLYGON 0 0 0.65 0 0.65 0.8 0 0.8 ;
      LAYER M1 ;
        POLYGON 0.159 0.541 0.323 0.541 0.323 0.263 0.04 0.263 0.04 0.091 0.115 0.091 0.115 0.202 0.373 0.202 0.373 0.375 0.458 0.375 0.458 0.425 0.373 0.425 0.373 0.592 0.231 0.592 0.231 0.709 0.159 0.709  ;
        POLYGON 0 -0.033 0.65 -0.033 0.65 0.033 0.621 0.033 0.621 0.161 0.549 0.161 0.549 0.033 0.361 0.033 0.361 0.127 0.289 0.127 0.289 0.033 0 0.033  ;
        POLYGON 0 0.767 0.029 0.767 0.029 0.545 0.101 0.545 0.101 0.767 0.289 0.767 0.289 0.656 0.361 0.656 0.361 0.767 0.549 0.767 0.549 0.639 0.621 0.639 0.621 0.767 0.65 0.767 0.65 0.833 0 0.833  ;
  END
END ISO_FENCE0N_X2_RVT_30

MACRO ISO_FENCE0N_X4_RVT_30
  CLASS core ;
  FOREIGN ISO_FENCE0N_X4_RVT_30 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CellTemplate ;
  SIZE 1.17 BY 0.8 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.03096 ;
    PORT
      LAYER M1 ;
        POLYGON 0.167 0.183 0.357 0.183 0.357 0.452 0.291 0.452 0.291 0.233 0.167 0.233  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.03096 ;
    PORT
      LAYER M2 ;
        POLYGON 0.077 0.425 0.588 0.425 0.588 0.475 0.077 0.475  ;
      LAYER V1 ;
        POLYGON 0.109 0.425 0.159 0.425 0.159 0.475 0.109 0.475  ;
        POLYGON 0.468 0.425 0.518 0.425 0.518 0.475 0.468 0.475  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.1032 ;
    PORT
      LAYER M1 ;
        POLYGON 0.679 0.54 0.945 0.54 0.945 0.258 0.679 0.258 0.679 0.091 0.751 0.091 0.751 0.208 0.939 0.208 0.939 0.091 1.011 0.091 1.011 0.709 0.939 0.709 0.939 0.59 0.751 0.59 0.751 0.709 0.679 0.709  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 0.735 1.17 0.735 1.17 0.865 0 0.865  ;
      LAYER V1 ;
        POLYGON 0.04 0.775 0.09 0.775 0.09 0.825 0.04 0.825  ;
        POLYGON 0.17 0.775 0.22 0.775 0.22 0.825 0.17 0.825  ;
        POLYGON 0.3 0.775 0.35 0.775 0.35 0.825 0.3 0.825  ;
        POLYGON 0.43 0.775 0.48 0.775 0.48 0.825 0.43 0.825  ;
        POLYGON 0.56 0.775 0.61 0.775 0.61 0.825 0.56 0.825  ;
        POLYGON 0.69 0.775 0.74 0.775 0.74 0.825 0.69 0.825  ;
        POLYGON 0.82 0.775 0.87 0.775 0.87 0.825 0.82 0.825  ;
        POLYGON 0.95 0.775 1 0.775 1 0.825 0.95 0.825  ;
        POLYGON 1.08 0.775 1.13 0.775 1.13 0.825 1.08 0.825  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 -0.065 1.17 -0.065 1.17 0.065 0 0.065  ;
      LAYER V1 ;
        POLYGON 0.04 -0.025 0.09 -0.025 0.09 0.025 0.04 0.025  ;
        POLYGON 0.17 -0.025 0.22 -0.025 0.22 0.025 0.17 0.025  ;
        POLYGON 0.3 -0.025 0.35 -0.025 0.35 0.025 0.3 0.025  ;
        POLYGON 0.43 -0.025 0.48 -0.025 0.48 0.025 0.43 0.025  ;
        POLYGON 0.56 -0.025 0.61 -0.025 0.61 0.025 0.56 0.025  ;
        POLYGON 0.69 -0.025 0.74 -0.025 0.74 0.025 0.69 0.025  ;
        POLYGON 0.82 -0.025 0.87 -0.025 0.87 0.025 0.82 0.025  ;
        POLYGON 0.95 -0.025 1 -0.025 1 0.025 0.95 0.025  ;
        POLYGON 1.08 -0.025 1.13 -0.025 1.13 0.025 1.08 0.025  ;
    END
  END VSS
  OBS
      LAYER RVT ;
        POLYGON 0 0 1.17 0 1.17 0.8 0 0.8 ;
      LAYER M1 ;
        POLYGON 0.159 0.543 0.578 0.543 0.578 0.252 0.446 0.252 0.446 0.133 0.161 0.133 0.161 0.083 0.499 0.083 0.499 0.202 0.628 0.202 0.628 0.375 0.713 0.375 0.713 0.425 0.628 0.425 0.628 0.593 0.491 0.593 0.491 0.709 0.419 0.709 0.419 0.593 0.231 0.593 0.231 0.709 0.159 0.709  ;
        POLYGON 0.095 0.292 0.167 0.292 0.167 0.485 0.095 0.485  ;
        POLYGON 0.454 0.31 0.526 0.31 0.526 0.485 0.454 0.485  ;
        POLYGON 0 -0.033 1.17 -0.033 1.17 0.033 1.141 0.033 1.141 0.223 1.069 0.223 1.069 0.033 0.881 0.033 0.881 0.144 0.809 0.144 0.809 0.033 0.621 0.033 0.621 0.144 0.549 0.144 0.549 0.033 0.101 0.033 0.101 0.224 0.029 0.224 0.029 0.033 0 0.033  ;
        POLYGON 0 0.767 0.029 0.767 0.029 0.565 0.101 0.565 0.101 0.767 0.289 0.767 0.289 0.656 0.361 0.656 0.361 0.767 0.549 0.767 0.549 0.656 0.621 0.656 0.621 0.767 0.809 0.767 0.809 0.656 0.881 0.656 0.881 0.767 1.069 0.767 1.069 0.577 1.141 0.577 1.141 0.767 1.17 0.767 1.17 0.833 0 0.833  ;
  END
END ISO_FENCE0N_X4_RVT_30

MACRO ISO_FENCE0_X1_RVT_30
  CLASS core ;
  FOREIGN ISO_FENCE0_X1_RVT_30 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X ;
  SITE CellTemplate ;
  SIZE 0.39 BY 0.8 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.01392 ;
    PORT
      LAYER M1 ;
        POLYGON 0.184 0.348 0.265 0.348 0.265 0.452 0.25 0.452 0.25 0.587 0.184 0.587  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.01392 ;
    PORT
      LAYER M1 ;
        POLYGON 0.059 0.348 0.134 0.348 0.134 0.452 0.125 0.452 0.125 0.584 0.059 0.584  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.040724 ;
    PORT
      LAYER M1 ;
        POLYGON 0.26 0.651 0.3 0.651 0.3 0.488 0.315 0.488 0.315 0.258 0.159 0.258 0.159 0.091 0.231 0.091 0.231 0.208 0.365 0.208 0.365 0.717 0.26 0.717  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 0.735 0.39 0.735 0.39 0.865 0 0.865  ;
      LAYER V1 ;
        POLYGON 0.04 0.775 0.09 0.775 0.09 0.825 0.04 0.825  ;
        POLYGON 0.17 0.775 0.22 0.775 0.22 0.825 0.17 0.825  ;
        POLYGON 0.3 0.775 0.35 0.775 0.35 0.825 0.3 0.825  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 -0.065 0.39 -0.065 0.39 0.065 0 0.065  ;
      LAYER V1 ;
        POLYGON 0.04 -0.025 0.09 -0.025 0.09 0.025 0.04 0.025  ;
        POLYGON 0.17 -0.025 0.22 -0.025 0.22 0.025 0.17 0.025  ;
        POLYGON 0.3 -0.025 0.35 -0.025 0.35 0.025 0.3 0.025  ;
    END
  END VSS
  OBS
      LAYER RVT ;
        POLYGON 0 0 0.39 0 0.39 0.8 0 0.8 ;
      LAYER M1 ;
        POLYGON 0 -0.033 0.39 -0.033 0.39 0.033 0.361 0.033 0.361 0.15 0.289 0.15 0.289 0.033 0.101 0.033 0.101 0.223 0.029 0.223 0.029 0.033 0 0.033  ;
        POLYGON 0 0.767 0.029 0.767 0.029 0.646 0.101 0.646 0.101 0.767 0.39 0.767 0.39 0.833 0 0.833  ;
  END
END ISO_FENCE0_X1_RVT_30

MACRO ISO_FENCE0_X2_RVT_30
  CLASS core ;
  FOREIGN ISO_FENCE0_X2_RVT_30 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CellTemplate ;
  SIZE 0.65 BY 0.8 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.02784 ;
    PORT
      LAYER M1 ;
        POLYGON 0.177 0.508 0.219 0.508 0.219 0.395 0.335 0.395 0.335 0.445 0.276 0.445 0.276 0.558 0.227 0.558 0.227 0.707 0.177 0.707  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.02784 ;
    PORT
      LAYER M1 ;
        POLYGON 0.055 0.368 0.11 0.368 0.11 0.295 0.499 0.295 0.499 0.348 0.525 0.348 0.525 0.452 0.449 0.452 0.449 0.345 0.169 0.345 0.169 0.434 0.127 0.434 0.127 0.517 0.055 0.517  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.067 ;
    PORT
      LAYER M1 ;
        POLYGON 0.289 0.622 0.419 0.622 0.419 0.543 0.575 0.543 0.575 0.245 0.159 0.245 0.159 0.187 0.625 0.187 0.625 0.593 0.485 0.593 0.485 0.678 0.361 0.678 0.361 0.717 0.289 0.717  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 0.735 0.65 0.735 0.65 0.865 0 0.865  ;
      LAYER V1 ;
        POLYGON 0.04 0.775 0.09 0.775 0.09 0.825 0.04 0.825  ;
        POLYGON 0.17 0.775 0.22 0.775 0.22 0.825 0.17 0.825  ;
        POLYGON 0.3 0.775 0.35 0.775 0.35 0.825 0.3 0.825  ;
        POLYGON 0.43 0.775 0.48 0.775 0.48 0.825 0.43 0.825  ;
        POLYGON 0.56 0.775 0.61 0.775 0.61 0.825 0.56 0.825  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 -0.065 0.65 -0.065 0.65 0.065 0 0.065  ;
      LAYER V1 ;
        POLYGON 0.04 -0.025 0.09 -0.025 0.09 0.025 0.04 0.025  ;
        POLYGON 0.17 -0.025 0.22 -0.025 0.22 0.025 0.17 0.025  ;
        POLYGON 0.3 -0.025 0.35 -0.025 0.35 0.025 0.3 0.025  ;
        POLYGON 0.43 -0.025 0.48 -0.025 0.48 0.025 0.43 0.025  ;
        POLYGON 0.56 -0.025 0.61 -0.025 0.61 0.025 0.56 0.025  ;
    END
  END VSS
  OBS
      LAYER RVT ;
        POLYGON 0 0 0.65 0 0.65 0.8 0 0.8 ;
      LAYER M1 ;
        POLYGON 0.421 0.087 0.549 0.087 0.549 0.033 0.361 0.033 0.361 0.125 0.289 0.125 0.289 0.033 0.101 0.033 0.101 0.237 0.029 0.237 0.029 0.033 0 0.033 0 -0.033 0.65 -0.033 0.65 0.033 0.621 0.033 0.621 0.137 0.421 0.137  ;
        POLYGON 0 0.767 0.029 0.767 0.029 0.581 0.101 0.581 0.101 0.767 0.549 0.767 0.549 0.651 0.621 0.651 0.621 0.767 0.65 0.767 0.65 0.833 0 0.833  ;
  END
END ISO_FENCE0_X2_RVT_30

MACRO ISO_FENCE0_X4_RVT_30
  CLASS core ;
  FOREIGN ISO_FENCE0_X4_RVT_30 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CellTemplate ;
  SIZE 1.17 BY 0.8 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.05568 ;
    PORT
      LAYER M1 ;
        POLYGON 0.284 0.395 0.454 0.395 0.454 0.464 0.729 0.464 0.729 0.395 0.883 0.395 0.883 0.464 0.779 0.464 0.779 0.514 0.388 0.514 0.388 0.464 0.284 0.464  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.05568 ;
    PORT
      LAYER M1 ;
        POLYGON 0.083 0.295 1.019 0.295 1.019 0.348 1.045 0.348 1.045 0.452 0.969 0.452 0.969 0.345 0.679 0.345 0.679 0.406 0.621 0.406 0.621 0.345 0.155 0.345 0.155 0.515 0.083 0.515  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.134 ;
    PORT
      LAYER M1 ;
        POLYGON 0.287 0.567 0.363 0.567 0.363 0.667 0.449 0.667 0.449 0.567 0.729 0.567 0.729 0.667 0.816 0.667 0.816 0.556 0.874 0.556 0.874 0.667 0.924 0.667 0.924 0.536 1.095 0.536 1.095 0.245 0.159 0.245 0.159 0.091 0.231 0.091 0.231 0.191 0.419 0.191 0.419 0.091 0.491 0.091 0.491 0.191 0.679 0.191 0.679 0.091 0.751 0.091 0.751 0.191 0.939 0.191 0.939 0.091 1.011 0.091 1.011 0.195 1.145 0.195 1.145 0.586 0.974 0.586 0.974 0.717 0.679 0.717 0.679 0.617 0.499 0.617 0.499 0.717 0.287 0.717  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 0.735 1.17 0.735 1.17 0.865 0 0.865  ;
      LAYER V1 ;
        POLYGON 0.04 0.775 0.09 0.775 0.09 0.825 0.04 0.825  ;
        POLYGON 0.17 0.775 0.22 0.775 0.22 0.825 0.17 0.825  ;
        POLYGON 0.3 0.775 0.35 0.775 0.35 0.825 0.3 0.825  ;
        POLYGON 0.43 0.775 0.48 0.775 0.48 0.825 0.43 0.825  ;
        POLYGON 0.56 0.775 0.61 0.775 0.61 0.825 0.56 0.825  ;
        POLYGON 0.69 0.775 0.74 0.775 0.74 0.825 0.69 0.825  ;
        POLYGON 0.82 0.775 0.87 0.775 0.87 0.825 0.82 0.825  ;
        POLYGON 0.95 0.775 1 0.775 1 0.825 0.95 0.825  ;
        POLYGON 1.08 0.775 1.13 0.775 1.13 0.825 1.08 0.825  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 -0.065 1.17 -0.065 1.17 0.065 0 0.065  ;
      LAYER V1 ;
        POLYGON 0.04 -0.025 0.09 -0.025 0.09 0.025 0.04 0.025  ;
        POLYGON 0.17 -0.025 0.22 -0.025 0.22 0.025 0.17 0.025  ;
        POLYGON 0.3 -0.025 0.35 -0.025 0.35 0.025 0.3 0.025  ;
        POLYGON 0.43 -0.025 0.48 -0.025 0.48 0.025 0.43 0.025  ;
        POLYGON 0.56 -0.025 0.61 -0.025 0.61 0.025 0.56 0.025  ;
        POLYGON 0.69 -0.025 0.74 -0.025 0.74 0.025 0.69 0.025  ;
        POLYGON 0.82 -0.025 0.87 -0.025 0.87 0.025 0.82 0.025  ;
        POLYGON 0.95 -0.025 1 -0.025 1 0.025 0.95 0.025  ;
        POLYGON 1.08 -0.025 1.13 -0.025 1.13 0.025 1.08 0.025  ;
    END
  END VSS
  OBS
      LAYER RVT ;
        POLYGON 0 0 1.17 0 1.17 0.8 0 0.8 ;
      LAYER M1 ;
        POLYGON 0 -0.033 1.17 -0.033 1.17 0.033 1.141 0.033 1.141 0.137 1.069 0.137 1.069 0.033 0.881 0.033 0.881 0.133 0.809 0.133 0.809 0.033 0.621 0.033 0.621 0.133 0.549 0.133 0.549 0.033 0.361 0.033 0.361 0.133 0.289 0.133 0.289 0.033 0.101 0.033 0.101 0.237 0.029 0.237 0.029 0.033 0 0.033  ;
        POLYGON 0 0.767 0.029 0.767 0.029 0.58 0.101 0.58 0.101 0.767 0.549 0.767 0.549 0.675 0.621 0.675 0.621 0.767 1.069 0.767 1.069 0.644 1.141 0.644 1.141 0.767 1.17 0.767 1.17 0.833 0 0.833  ;
  END
END ISO_FENCE0_X4_RVT_30

MACRO ISO_FENCE1N_X1_RVT_30
  CLASS core ;
  FOREIGN ISO_FENCE1N_X1_RVT_30 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X ;
  SITE CellTemplate ;
  SIZE 0.39 BY 0.8 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.0147 ;
    PORT
      LAYER M1 ;
        POLYGON 0.193 0.213 0.249 0.213 0.249 0.348 0.265 0.348 0.265 0.452 0.193 0.452  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.01509 ;
    PORT
      LAYER M1 ;
        POLYGON 0.071 0.291 0.143 0.291 0.143 0.498 0.071 0.498  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.04361 ;
    PORT
      LAYER M1 ;
        POLYGON 0.159 0.555 0.315 0.555 0.315 0.276 0.3 0.276 0.3 0.141 0.251 0.141 0.251 0.083 0.365 0.083 0.365 0.613 0.159 0.613  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 0.735 0.39 0.735 0.39 0.865 0 0.865  ;
      LAYER V1 ;
        POLYGON 0.04 0.775 0.09 0.775 0.09 0.825 0.04 0.825  ;
        POLYGON 0.17 0.775 0.22 0.775 0.22 0.825 0.17 0.825  ;
        POLYGON 0.3 0.775 0.35 0.775 0.35 0.825 0.3 0.825  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 -0.065 0.39 -0.065 0.39 0.065 0 0.065  ;
      LAYER V1 ;
        POLYGON 0.04 -0.025 0.09 -0.025 0.09 0.025 0.04 0.025  ;
        POLYGON 0.17 -0.025 0.22 -0.025 0.22 0.025 0.17 0.025  ;
        POLYGON 0.3 -0.025 0.35 -0.025 0.35 0.025 0.3 0.025  ;
    END
  END VSS
  OBS
      LAYER RVT ;
        POLYGON 0 0 0.39 0 0.39 0.8 0 0.8 ;
      LAYER M1 ;
        POLYGON 0 -0.033 0.39 -0.033 0.39 0.033 0.101 0.033 0.101 0.216 0.029 0.216 0.029 0.033 0 0.033  ;
        POLYGON 0 0.767 0.029 0.767 0.029 0.584 0.101 0.584 0.101 0.767 0.289 0.767 0.289 0.713 0.2 0.713 0.2 0.663 0.361 0.663 0.361 0.767 0.39 0.767 0.39 0.833 0 0.833  ;
  END
END ISO_FENCE1N_X1_RVT_30

MACRO ISO_FENCE1N_X2_RVT_30
  CLASS core ;
  FOREIGN ISO_FENCE1N_X2_RVT_30 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CellTemplate ;
  SIZE 0.65 BY 0.8 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.0294 ;
    PORT
      LAYER M1 ;
        POLYGON 0.173 0.091 0.239 0.091 0.239 0.282 0.255 0.282 0.255 0.354 0.359 0.354 0.359 0.405 0.205 0.405 0.205 0.332 0.189 0.332 0.189 0.21 0.173 0.21  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.03018 ;
    PORT
      LAYER M1 ;
        POLYGON 0.08 0.377 0.155 0.377 0.155 0.455 0.449 0.455 0.449 0.348 0.525 0.348 0.525 0.452 0.499 0.452 0.499 0.505 0.08 0.505  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.0735 ;
    PORT
      LAYER M1 ;
        POLYGON 0.159 0.555 0.575 0.555 0.575 0.245 0.289 0.245 0.289 0.091 0.361 0.091 0.361 0.195 0.625 0.195 0.625 0.613 0.159 0.613  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 0.735 0.65 0.735 0.65 0.865 0 0.865  ;
      LAYER V1 ;
        POLYGON 0.04 0.775 0.09 0.775 0.09 0.825 0.04 0.825  ;
        POLYGON 0.17 0.775 0.22 0.775 0.22 0.825 0.17 0.825  ;
        POLYGON 0.3 0.775 0.35 0.775 0.35 0.825 0.3 0.825  ;
        POLYGON 0.43 0.775 0.48 0.775 0.48 0.825 0.43 0.825  ;
        POLYGON 0.56 0.775 0.61 0.775 0.61 0.825 0.56 0.825  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 -0.065 0.65 -0.065 0.65 0.065 0 0.065  ;
      LAYER V1 ;
        POLYGON 0.04 -0.025 0.09 -0.025 0.09 0.025 0.04 0.025  ;
        POLYGON 0.17 -0.025 0.22 -0.025 0.22 0.025 0.17 0.025  ;
        POLYGON 0.3 -0.025 0.35 -0.025 0.35 0.025 0.3 0.025  ;
        POLYGON 0.43 -0.025 0.48 -0.025 0.48 0.025 0.43 0.025  ;
        POLYGON 0.56 -0.025 0.61 -0.025 0.61 0.025 0.56 0.025  ;
    END
  END VSS
  OBS
      LAYER RVT ;
        POLYGON 0 0 0.65 0 0.65 0.8 0 0.8 ;
      LAYER M1 ;
        POLYGON 0 -0.033 0.65 -0.033 0.65 0.033 0.621 0.033 0.621 0.137 0.549 0.137 0.549 0.033 0.101 0.033 0.101 0.298 0.029 0.298 0.029 0.033 0 0.033  ;
        POLYGON 0 0.767 0.029 0.767 0.029 0.563 0.101 0.563 0.101 0.767 0.289 0.767 0.289 0.675 0.361 0.675 0.361 0.767 0.549 0.767 0.549 0.713 0.421 0.713 0.421 0.663 0.621 0.663 0.621 0.767 0.65 0.767 0.65 0.833 0 0.833  ;
  END
END ISO_FENCE1N_X2_RVT_30

MACRO ISO_FENCE1N_X4_RVT_30
  CLASS core ;
  FOREIGN ISO_FENCE1N_X4_RVT_30 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CellTemplate ;
  SIZE 1.17 BY 0.8 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.0588 ;
    PORT
      LAYER M1 ;
        POLYGON 0.213 0.333 0.329 0.333 0.329 0.193 0.379 0.193 0.379 0.283 0.816 0.283 0.816 0.333 0.884 0.333 0.884 0.405 0.744 0.405 0.744 0.333 0.426 0.333 0.426 0.405 0.213 0.405  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.06036 ;
    PORT
      LAYER M1 ;
        POLYGON 0.089 0.302 0.155 0.302 0.155 0.455 0.479 0.455 0.479 0.383 0.694 0.383 0.694 0.455 0.969 0.455 0.969 0.348 1.045 0.348 1.045 0.452 1.019 0.452 1.019 0.505 0.644 0.505 0.644 0.444 0.529 0.444 0.529 0.505 0.089 0.505  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.147 ;
    PORT
      LAYER M1 ;
        POLYGON 0.159 0.555 1.095 0.555 1.095 0.258 0.89 0.258 0.89 0.133 0.744 0.133 0.744 0.233 0.429 0.233 0.429 0.133 0.161 0.133 0.161 0.083 0.479 0.083 0.479 0.183 0.694 0.183 0.694 0.083 0.94 0.083 0.94 0.208 1.145 0.208 1.145 0.605 1.011 0.605 1.011 0.709 0.939 0.709 0.939 0.609 0.751 0.609 0.751 0.709 0.679 0.709 0.679 0.609 0.491 0.609 0.491 0.709 0.419 0.709 0.419 0.609 0.231 0.609 0.231 0.709 0.159 0.709  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 0.735 1.17 0.735 1.17 0.865 0 0.865  ;
      LAYER V1 ;
        POLYGON 0.04 0.775 0.09 0.775 0.09 0.825 0.04 0.825  ;
        POLYGON 0.17 0.775 0.22 0.775 0.22 0.825 0.17 0.825  ;
        POLYGON 0.3 0.775 0.35 0.775 0.35 0.825 0.3 0.825  ;
        POLYGON 0.43 0.775 0.48 0.775 0.48 0.825 0.43 0.825  ;
        POLYGON 0.56 0.775 0.61 0.775 0.61 0.825 0.56 0.825  ;
        POLYGON 0.69 0.775 0.74 0.775 0.74 0.825 0.69 0.825  ;
        POLYGON 0.82 0.775 0.87 0.775 0.87 0.825 0.82 0.825  ;
        POLYGON 0.95 0.775 1 0.775 1 0.825 0.95 0.825  ;
        POLYGON 1.08 0.775 1.13 0.775 1.13 0.825 1.08 0.825  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 -0.065 1.17 -0.065 1.17 0.065 0 0.065  ;
      LAYER V1 ;
        POLYGON 0.04 -0.025 0.09 -0.025 0.09 0.025 0.04 0.025  ;
        POLYGON 0.17 -0.025 0.22 -0.025 0.22 0.025 0.17 0.025  ;
        POLYGON 0.3 -0.025 0.35 -0.025 0.35 0.025 0.3 0.025  ;
        POLYGON 0.43 -0.025 0.48 -0.025 0.48 0.025 0.43 0.025  ;
        POLYGON 0.56 -0.025 0.61 -0.025 0.61 0.025 0.56 0.025  ;
        POLYGON 0.69 -0.025 0.74 -0.025 0.74 0.025 0.69 0.025  ;
        POLYGON 0.82 -0.025 0.87 -0.025 0.87 0.025 0.82 0.025  ;
        POLYGON 0.95 -0.025 1 -0.025 1 0.025 0.95 0.025  ;
        POLYGON 1.08 -0.025 1.13 -0.025 1.13 0.025 1.08 0.025  ;
    END
  END VSS
  OBS
      LAYER RVT ;
        POLYGON 0 0 1.17 0 1.17 0.8 0 0.8 ;
      LAYER M1 ;
        POLYGON 0 -0.033 1.17 -0.033 1.17 0.033 1.141 0.033 1.141 0.15 1.069 0.15 1.069 0.033 0.621 0.033 0.621 0.125 0.549 0.125 0.549 0.033 0.101 0.033 0.101 0.24 0.029 0.24 0.029 0.033 0 0.033  ;
        POLYGON 0 0.767 0.029 0.767 0.029 0.563 0.101 0.563 0.101 0.767 0.289 0.767 0.289 0.667 0.361 0.667 0.361 0.767 0.549 0.767 0.549 0.667 0.621 0.667 0.621 0.767 0.809 0.767 0.809 0.667 0.881 0.667 0.881 0.767 1.069 0.767 1.069 0.663 1.141 0.663 1.141 0.767 1.17 0.767 1.17 0.833 0 0.833  ;
  END
END ISO_FENCE1N_X4_RVT_30

MACRO ISO_FENCE1_X1_RVT_30
  CLASS core ;
  FOREIGN ISO_FENCE1_X1_RVT_30 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CellTemplate ;
  SIZE 0.52 BY 0.8 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.00774 ;
    PORT
      LAYER M1 ;
        POLYGON 0.083 0.313 0.155 0.313 0.155 0.465 0.083 0.465  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.00774 ;
    PORT
      LAYER M1 ;
        POLYGON 0.207 0.313 0.273 0.313 0.273 0.465 0.207 0.465  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.040248 ;
    PORT
      LAYER M1 ;
        POLYGON 0.419 0.612 0.43 0.612 0.43 0.488 0.445 0.488 0.445 0.301 0.43 0.301 0.43 0.166 0.411 0.166 0.411 0.091 0.495 0.091 0.495 0.709 0.419 0.709  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 0.735 0.52 0.735 0.52 0.865 0 0.865  ;
      LAYER V1 ;
        POLYGON 0.04 0.775 0.09 0.775 0.09 0.825 0.04 0.825  ;
        POLYGON 0.17 0.775 0.22 0.775 0.22 0.825 0.17 0.825  ;
        POLYGON 0.3 0.775 0.35 0.775 0.35 0.825 0.3 0.825  ;
        POLYGON 0.43 0.775 0.48 0.775 0.48 0.825 0.43 0.825  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 -0.065 0.52 -0.065 0.52 0.065 0 0.065  ;
      LAYER V1 ;
        POLYGON 0.04 -0.025 0.09 -0.025 0.09 0.025 0.04 0.025  ;
        POLYGON 0.17 -0.025 0.22 -0.025 0.22 0.025 0.17 0.025  ;
        POLYGON 0.3 -0.025 0.35 -0.025 0.35 0.025 0.3 0.025  ;
        POLYGON 0.43 -0.025 0.48 -0.025 0.48 0.025 0.43 0.025  ;
    END
  END VSS
  OBS
      LAYER RVT ;
        POLYGON 0 0 0.52 0 0.52 0.8 0 0.8 ;
      LAYER M1 ;
        POLYGON 0.04 0.523 0.323 0.523 0.323 0.252 0.159 0.252 0.159 0.091 0.231 0.091 0.231 0.202 0.373 0.202 0.373 0.348 0.395 0.348 0.395 0.452 0.373 0.452 0.373 0.576 0.115 0.576 0.115 0.709 0.04 0.709  ;
        POLYGON 0 -0.033 0.52 -0.033 0.52 0.033 0.361 0.033 0.361 0.144 0.289 0.144 0.289 0.033 0.101 0.033 0.101 0.248 0.029 0.248 0.029 0.033 0 0.033  ;
        POLYGON 0 0.767 0.289 0.767 0.289 0.656 0.361 0.656 0.361 0.767 0.52 0.767 0.52 0.833 0 0.833  ;
  END
END ISO_FENCE1_X1_RVT_30

MACRO ISO_FENCE1_X2_RVT_30
  CLASS core ;
  FOREIGN ISO_FENCE1_X2_RVT_30 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CellTemplate ;
  SIZE 0.65 BY 0.8 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.01548 ;
    PORT
      LAYER M1 ;
        POLYGON 0.083 0.316 0.155 0.316 0.155 0.468 0.083 0.468  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.01548 ;
    PORT
      LAYER M1 ;
        POLYGON 0.207 0.316 0.273 0.316 0.273 0.468 0.207 0.468  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.0516 ;
    PORT
      LAYER M1 ;
        POLYGON 0.423 0.471 0.556 0.471 0.556 0.289 0.423 0.289 0.423 0.091 0.489 0.091 0.489 0.235 0.606 0.235 0.606 0.521 0.489 0.521 0.489 0.709 0.423 0.709  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 0.735 0.65 0.735 0.65 0.865 0 0.865  ;
      LAYER V1 ;
        POLYGON 0.04 0.775 0.09 0.775 0.09 0.825 0.04 0.825  ;
        POLYGON 0.17 0.775 0.22 0.775 0.22 0.825 0.17 0.825  ;
        POLYGON 0.3 0.775 0.35 0.775 0.35 0.825 0.3 0.825  ;
        POLYGON 0.43 0.775 0.48 0.775 0.48 0.825 0.43 0.825  ;
        POLYGON 0.56 0.775 0.61 0.775 0.61 0.825 0.56 0.825  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 -0.065 0.65 -0.065 0.65 0.065 0 0.065  ;
      LAYER V1 ;
        POLYGON 0.04 -0.025 0.09 -0.025 0.09 0.025 0.04 0.025  ;
        POLYGON 0.17 -0.025 0.22 -0.025 0.22 0.025 0.17 0.025  ;
        POLYGON 0.3 -0.025 0.35 -0.025 0.35 0.025 0.3 0.025  ;
        POLYGON 0.43 -0.025 0.48 -0.025 0.48 0.025 0.43 0.025  ;
        POLYGON 0.56 -0.025 0.61 -0.025 0.61 0.025 0.56 0.025  ;
    END
  END VSS
  OBS
      LAYER RVT ;
        POLYGON 0 0 0.65 0 0.65 0.8 0 0.8 ;
      LAYER M1 ;
        POLYGON 0.04 0.526 0.323 0.526 0.323 0.258 0.159 0.258 0.159 0.091 0.231 0.091 0.231 0.208 0.373 0.208 0.373 0.371 0.459 0.371 0.459 0.421 0.373 0.421 0.373 0.576 0.115 0.576 0.115 0.709 0.04 0.709  ;
        POLYGON 0 -0.033 0.65 -0.033 0.65 0.033 0.621 0.033 0.621 0.177 0.549 0.177 0.549 0.033 0.361 0.033 0.361 0.144 0.289 0.144 0.289 0.033 0.101 0.033 0.101 0.254 0.029 0.254 0.029 0.033 0 0.033  ;
        POLYGON 0 0.767 0.289 0.767 0.289 0.656 0.361 0.656 0.361 0.767 0.549 0.767 0.549 0.579 0.621 0.579 0.621 0.767 0.65 0.767 0.65 0.833 0 0.833  ;
  END
END ISO_FENCE1_X2_RVT_30

MACRO ISO_FENCE1_X4_RVT_30
  CLASS core ;
  FOREIGN ISO_FENCE1_X4_RVT_30 0.0 0.0 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y ;
  SITE CellTemplate ;
  SIZE 1.17 BY 0.8 ;
  PIN A
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.03096 ;
    PORT
      LAYER M1 ;
        POLYGON 0.21 0.536 0.3 0.536 0.3 0.313 0.366 0.313 0.366 0.586 0.21 0.586  ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    ANTENNAGATEAREA 0.03096 ;
    PORT
      LAYER M2 ;
        POLYGON 0.077 0.325 0.542 0.325 0.542 0.375 0.077 0.375  ;
      LAYER V1 ;
        POLYGON 0.109 0.325 0.159 0.325 0.159 0.375 0.109 0.375  ;
        POLYGON 0.46 0.325 0.51 0.325 0.51 0.375 0.46 0.375  ;
    END
  END EN
  PIN Z
    DIRECTION OUTPUT ;
    ANTENNADIFFAREA 0.1032 ;
    PORT
      LAYER M1 ;
        POLYGON 0.679 0.471 0.95 0.471 0.95 0.283 0.679 0.283 0.679 0.091 0.751 0.091 0.751 0.233 0.939 0.233 0.939 0.091 1.011 0.091 1.011 0.709 0.939 0.709 0.939 0.521 0.751 0.521 0.751 0.709 0.679 0.709  ;
    END
  END Z
  PIN VDD
    DIRECTION INOUT ;
    USE power ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 0.735 1.17 0.735 1.17 0.865 0 0.865  ;
      LAYER V1 ;
        POLYGON 0.04 0.775 0.09 0.775 0.09 0.825 0.04 0.825  ;
        POLYGON 0.17 0.775 0.22 0.775 0.22 0.825 0.17 0.825  ;
        POLYGON 0.3 0.775 0.35 0.775 0.35 0.825 0.3 0.825  ;
        POLYGON 0.43 0.775 0.48 0.775 0.48 0.825 0.43 0.825  ;
        POLYGON 0.56 0.775 0.61 0.775 0.61 0.825 0.56 0.825  ;
        POLYGON 0.69 0.775 0.74 0.775 0.74 0.825 0.69 0.825  ;
        POLYGON 0.82 0.775 0.87 0.775 0.87 0.825 0.82 0.825  ;
        POLYGON 0.95 0.775 1 0.775 1 0.825 0.95 0.825  ;
        POLYGON 1.08 0.775 1.13 0.775 1.13 0.825 1.08 0.825  ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE ground ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        POLYGON 0 -0.065 1.17 -0.065 1.17 0.065 0 0.065  ;
      LAYER V1 ;
        POLYGON 0.04 -0.025 0.09 -0.025 0.09 0.025 0.04 0.025  ;
        POLYGON 0.17 -0.025 0.22 -0.025 0.22 0.025 0.17 0.025  ;
        POLYGON 0.3 -0.025 0.35 -0.025 0.35 0.025 0.3 0.025  ;
        POLYGON 0.43 -0.025 0.48 -0.025 0.48 0.025 0.43 0.025  ;
        POLYGON 0.56 -0.025 0.61 -0.025 0.61 0.025 0.56 0.025  ;
        POLYGON 0.69 -0.025 0.74 -0.025 0.74 0.025 0.69 0.025  ;
        POLYGON 0.82 -0.025 0.87 -0.025 0.87 0.025 0.82 0.025  ;
        POLYGON 0.95 -0.025 1 -0.025 1 0.025 0.95 0.025  ;
        POLYGON 1.08 -0.025 1.13 -0.025 1.13 0.025 1.08 0.025  ;
    END
  END VSS
  OBS
      LAYER RVT ;
        POLYGON 0 0 1.17 0 1.17 0.8 0 0.8 ;
      LAYER M1 ;
        POLYGON 0.161 0.667 0.444 0.667 0.444 0.548 0.576 0.548 0.576 0.248 0.159 0.248 0.159 0.091 0.231 0.091 0.231 0.183 0.626 0.183 0.626 0.363 0.892 0.363 0.892 0.421 0.626 0.421 0.626 0.598 0.497 0.598 0.497 0.717 0.161 0.717  ;
        POLYGON 0.09 0.306 0.162 0.306 0.162 0.467 0.09 0.467  ;
        POLYGON 0.46 0.308 0.526 0.308 0.526 0.464 0.46 0.464  ;
        POLYGON 0 -0.033 1.17 -0.033 1.17 0.033 1.141 0.033 1.141 0.26 1.069 0.26 1.069 0.033 0.881 0.033 0.881 0.144 0.809 0.144 0.809 0.033 0.621 0.033 0.621 0.125 0.549 0.125 0.549 0.033 0.361 0.033 0.361 0.125 0.289 0.125 0.289 0.033 0.101 0.033 0.101 0.229 0.029 0.229 0.029 0.033 0 0.033  ;
        POLYGON 0 0.767 0.029 0.767 0.029 0.563 0.101 0.563 0.101 0.767 0.549 0.767 0.549 0.656 0.621 0.656 0.621 0.767 0.809 0.767 0.809 0.579 0.881 0.579 0.881 0.767 1.069 0.767 1.069 0.467 1.141 0.467 1.141 0.767 1.17 0.767 1.17 0.833 0 0.833  ;
  END
END ISO_FENCE1_X4_RVT_30

END LIBRARY
#
# End of file
#
